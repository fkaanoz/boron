
module dec_key_scheduler();



endmodule
