`timescale 1ns/1ps


module round_permutation();


endmodule
