
module encrytion();



endmodule
