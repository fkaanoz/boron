
module dec_sbox_bank();


endmodule
