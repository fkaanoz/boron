`timescale 1ns/1ps


module dec_round_permutation();


endmodule
