
module dec_xor_operation();


endmodule
