
module dec_sbox_layer();


endmodule
