
module dec_sbox();


endmodule
