`timescale 1ns/1ps


module boron(
    input clk,
    input reset,
    input [63:0] plain_text,
    input [79:0] master_key

    output enc_done,
    output [63:0] cipher_text

);



endmodule
