`timescale 1ns/1ps


module dec_sbox_bank();


endmodule
