`timescale 1ns/1ps


module sbox_layer();


endmodule
