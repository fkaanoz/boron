`timescale 1ns/1ps


module dec_key_scheduler();



endmodule
