
module dec_block_shuffle();


endmodule
