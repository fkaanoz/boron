`timescale 1ns/1ps


module dec_xor_operation();


endmodule
