`timescale 1ns/1ps


module dec_sbox_layer();


endmodule
