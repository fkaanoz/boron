
module block_shuffle();


endmodule
