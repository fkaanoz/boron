`timescale 1ns/1ps


module decrytion();



endmodule
