
module sbox();


endmodule
