`timescale 1ns/1ps


module dec_block_shuffle();


endmodule
