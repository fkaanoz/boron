
module decrytion();



endmodule
