`timescale 1ns/1ps


module encrytion();



endmodule
