
module round_permutation();


endmodule
