`timescale 1ns/1ps


module enc_key_scheduler();


endmodule
