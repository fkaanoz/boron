
module sbox_layer();


endmodule
