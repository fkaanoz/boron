
module xor_operation();


endmodule
