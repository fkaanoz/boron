`timescale 1ns/1ps


module xor_operation();


endmodule
