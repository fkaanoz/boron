
module dec_round_permutation();


endmodule
