
module enc_key_scheduler();


endmodule
