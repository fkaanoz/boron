`timescale 1ns/1ps


module block_shuffle();


endmodule
