
module sbox_bank();


endmodule
