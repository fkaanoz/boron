`timescale 1ns/1ps


module sbox();


endmodule
